netcdf test {

dimensions:
	time = unlimited ; // (0 currently)
	X = 4 ;
	
variables:
	int A(time, X) ;
	    	A:_FillValue = -99 ;
	        A:att1 = "ASCII text attribute" ;
A:att2 = 3.14 ;
		A:att3 = 42 ;
		A:att4 = 1.1, 2, 0.5 ;
		A:att5 = 1, 2 ;
		A:att6 = 1.f, 2 ;
		A:att7 = 1.2f, 1.3e18, 1.0e21 ;
		A:att8 = 3s, 11 ;
		A:att9 = "Bjørn Ådlandsvik" ;
// Comment to separate global attributes
   	  :type = "Handwritten input for testing" ;
}


